module DebounceTest;


initial begin

    #5000;

    #50000;
    $finish;
    
end
endmodule